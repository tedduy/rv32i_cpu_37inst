// =============================================================================
// Sequence: TC 1.1.9 - OR Instruction
// =============================================================================
// Category: ISA Coverage
// Priority: CRITICAL
// Description: Bitwise OR
// =============================================================================

class tc_1_1_9_or_seq extends uvm_sequence #(rv32i_transaction);
    
    `uvm_object_utils(tc_1_1_9_or_seq)
    
    function new(string name = "tc_1_1_9_or_seq");
        super.new(name);
    endfunction
    
    task body();
        rv32i_transaction tr;
        
        `uvm_info(get_type_name(), "Starting OR sequence", UVM_MEDIUM)
        
        // ======================================================================
        // Test Case: OR - Bitwise OR
        // ======================================================================
        tr = rv32i_transaction::type_id::create("or_test");
        start_item(tr);
        
        tr.test_name = "OR Test";
        // TODO: Configure instruction encoding and test values
        // tr.opcode = ...;
        // tr.funct3 = ...;
        // tr.rd = ...;
        // tr.rs1 = ...;
        // tr.rs2 = ...;
        // tr.instruction = {tr.funct7, tr.rs2, tr.rs1, tr.funct3, tr.rd, tr.opcode};
        
        finish_item(tr);
        `uvm_info(get_type_name(), "Sent: OR test transaction", UVM_HIGH)
        
        `uvm_info(get_type_name(), "OR sequence completed", UVM_MEDIUM)
        
    endtask

endclass : tc_1_1_9_or_seq
