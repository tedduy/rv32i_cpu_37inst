// =============================================================================
// Sequence: TC 6.4.2 - STORE_LOAD_FORWARD Instruction
// =============================================================================
// Category: Memory System
// Priority: HIGH
// Description: Store-to-load forwarding
// =============================================================================

class tc_6_4_2_store_load_forward_seq extends uvm_sequence #(rv32i_transaction);
    
    `uvm_object_utils(tc_6_4_2_store_load_forward_seq)
    
    function new(string name = "tc_6_4_2_store_load_forward_seq");
        super.new(name);
    endfunction
    
    task body();
        rv32i_transaction tr;
        
        `uvm_info(get_type_name(), "Starting STORE_LOAD_FORWARD sequence", UVM_MEDIUM)
        
        // ======================================================================
        // Test Case: STORE_LOAD_FORWARD - Store-to-load forwarding
        // ======================================================================
        tr = rv32i_transaction::type_id::create("store_load_forward_test");
        start_item(tr);
        
        tr.test_name = "STORE_LOAD_FORWARD Test";
        // TODO: Configure instruction encoding and test values
        // tr.opcode = ...;
        // tr.funct3 = ...;
        // tr.rd = ...;
        // tr.rs1 = ...;
        // tr.rs2 = ...;
        // tr.instruction = {tr.funct7, tr.rs2, tr.rs1, tr.funct3, tr.rd, tr.opcode};
        
        finish_item(tr);
        `uvm_info(get_type_name(), "Sent: STORE_LOAD_FORWARD test transaction", UVM_HIGH)
        
        `uvm_info(get_type_name(), "STORE_LOAD_FORWARD sequence completed", UVM_MEDIUM)
        
    endtask

endclass : tc_6_4_2_store_load_forward_seq
