// =============================================================================
// Sequence: TC 9.3.1 - LOAD_FORWARD Instruction
// =============================================================================
// Category: Forwarding Paths
// Priority: CRITICAL
// Description: Load result forwarding
// =============================================================================

class tc_9_3_1_load_forward_seq extends uvm_sequence #(rv32i_transaction);
    
    `uvm_object_utils(tc_9_3_1_load_forward_seq)
    
    function new(string name = "tc_9_3_1_load_forward_seq");
        super.new(name);
    endfunction
    
    task body();
        rv32i_transaction tr;
        
        `uvm_info(get_type_name(), "Starting LOAD_FORWARD sequence", UVM_MEDIUM)
        
        // ======================================================================
        // Test Case: LOAD_FORWARD - Load result forwarding
        // ======================================================================
        tr = rv32i_transaction::type_id::create("load_forward_test");
        start_item(tr);
        
        tr.test_name = "LOAD_FORWARD Test";
        // TODO: Configure instruction encoding and test values
        // tr.opcode = ...;
        // tr.funct3 = ...;
        // tr.rd = ...;
        // tr.rs1 = ...;
        // tr.rs2 = ...;
        // tr.instruction = {tr.funct7, tr.rs2, tr.rs1, tr.funct3, tr.rd, tr.opcode};
        
        finish_item(tr);
        `uvm_info(get_type_name(), "Sent: LOAD_FORWARD test transaction", UVM_HIGH)
        
        `uvm_info(get_type_name(), "LOAD_FORWARD sequence completed", UVM_MEDIUM)
        
    endtask

endclass : tc_9_3_1_load_forward_seq
