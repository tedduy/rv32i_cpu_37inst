module Instruction_Mem #(
	parameter N = 32,
    parameter DEPTH = 76
)(
	input logic  i_clk,
    input logic  i_arst_n,		 // Reset active low	
  	input logic  [N-1:0] i_addr, // Address
  	output logic [N-1:0] o_inst  // Instruction
);
  //76 words, each word N bits
  logic [N-1:0] Imemory [0:DEPTH - 1];
  
  localparam int ADDR_LSB = 2;
  localparam int INDEX_W  = $clog2(DEPTH);
  wire [INDEX_W-1:0] word_idx = i_addr[ADDR_LSB +: INDEX_W];
  
  int i;
  
  assign o_inst = Imemory[word_idx];
   
  always_ff @(posedge i_clk or negedge i_arst_n) begin
    if(!i_arst_n) begin 
       for(i = 0; i < DEPTH; i = i + 1) begin
         Imemory[i] = '0;
       end

    end else begin
            Imemory[0]  = 32'b00000000000000000000000000000000; // 0x00000000 | nop (encoded as 0)

      // ===== R-type (rs1, rs2 ∈ {x1,x2,x4,x5}; rd ∈ {x3,x6}) =====
      Imemory[1]  = 32'b00000000001000001000000110110011; // 0x002081b3 | add x3, x1, x2
      Imemory[2]  = 32'b01000000010100100000011000110011; // 0x40520333 | sub x6, x4, x5
      Imemory[3]  = 32'b00000000010000001001000110110011; // 0x004091b3 | sll x3, x1, x4
      Imemory[4]  = 32'b00000000010100010010011000110011; // 0x00512333 | slt x6, x2, x5
      Imemory[5]  = 32'b00000000010000101011000110110011; // 0x0042b1b3 | sltu x3, x5, x4
      Imemory[6]  = 32'b00000000010100001100011000110011; // 0x0050c333 | xor x6, x1, x5
      Imemory[7]  = 32'b00000000001000100101000110110011; // 0x002251b3 | srl x3, x4, x2
      Imemory[8]  = 32'b01000000000100101101011000110011; // 0x4012d333 | sra x6, x5, x1
      Imemory[9]  = 32'b00000000010000001110000110110011; // 0x0040e1b3 | or  x3, x1, x4
      Imemory[10] = 32'b00000000010100010111011000110011; // 0x00517333 | and x6, x2, x5
      Imemory[11] = 32'b00000000010000101100011000110011; // 0x0042c333 | add x6, x5, x4
      Imemory[12] = 32'b01000000000100010000000110110011; // 0x401101b3 | sub x3, x2, x1
      Imemory[13] = 32'b00000000010000010001011000110011; // 0x004115b3 | sll x6, x2, x4
      Imemory[14] = 32'b00000000010100001010000110110011; // 0x0050a1b3 | slt x3, x1, x5
      Imemory[15] = 32'b00000000010100100110011000110011; // 0x00526633 | sltu x6, x4, x5
      Imemory[16] = 32'b00000000010000010100000110110011; // 0x004141b3 | xor x3, x2, x4
      Imemory[17] = 32'b00000000000100100101011000110011; // 0x001255b3 | srl x6, x4, x1
      Imemory[18] = 32'b01000000001000101101000110110011; // 0x4022d1b3 | sra x3, x5, x2
      Imemory[19] = 32'b00000000001000100110011000110011; // 0x00226633 | or  x6, x4, x2
      Imemory[20] = 32'b00000000010100001111000110110011; // 0x0050f1b3 | and x3, x1, x5

      // ===== I-type (giống R-type: rd ∈ {x3,x6}; rs1 ∈ {x1,x2,x4,x5}) =====
      Imemory[21] = 32'b00000000110000001000000110010011; // 0x000c0193 | addi  x3, x1, 100
      Imemory[22] = 32'b11111100111000010000011000010011; // 0xffc10613 | addi  x6, x2, -50
      Imemory[23] = 32'b00000001100100100010000110010011; // 0x01922193 | slti  x3, x4, 25
      Imemory[24] = 32'b11111110111000101010011000010011; // 0xffe2a613 | slti  x6, x5, -10
      Imemory[25] = 32'b00001100100000001011011000010011; // 0x0c801613 | sltiu x6, x1, 200
      Imemory[26] = 32'b00000000111100010011000110010011; // 0x00f13193 | sltiu x3, x2, 15
      Imemory[27] = 32'b00000000111100101100011000010011; // 0x00f2c613 | xori  x6, x5, 255
      Imemory[28] = 32'b00000000010100100100000110010011; // 0x00524193 | xori  x3, x4, 85
      Imemory[29] = 32'b00000000000000001110000110010011; // 0x0000e193 | ori   x3, x1, 15
      Imemory[30] = 32'b00000000100000010110011000010011; // 0x00817613 | ori   x6, x2, 128
      Imemory[31] = 32'b00000000111100011111011000010011; // 0x00f1f613 | andi  x6, x3, 240
      Imemory[32] = 32'b00000000111100110111100110010011; // 0x00f37f93 | andi  x3, x6, 255
      Imemory[33] = 32'b00000000001100001001000110010011; // 0x00309193 | slli  x3, x1, 3
      Imemory[34] = 32'b00000000100000010001011000010011; // 0x00811593 | slli  x6, x2, 8
      Imemory[35] = 32'b00000000010000101101000110010011; // 0x0042d193 | srli  x3, x5, 4
      Imemory[36] = 32'b00000000110000001101011000010011; // 0x00c0d613 | srli  x6, x1, 12
      Imemory[37] = 32'b01000000001000100101000110010011; // 0x40225193 | srai  x3, x4, 2
      Imemory[38] = 32'b01000000011000010101011000010011; // 0x40615513 | srai  x6, x2, 6
      Imemory[39] = 32'b11111111111100101111000110010011; // 0xfff2f193 | addi  x3, x5, -1

      // ===== LOADs (I-type, rd ∈ {x3,x6}; base rs1 ∈ {x1,x2,x4,x5}) =====
      Imemory[40] = 32'b00000000101000010000000110000011; // 0x00a10183 | lb   x3, 10(x2)
      Imemory[41] = 32'b11111111001100000000011000000011; // 0xff300603 | lb   x6, -5(x1)
      Imemory[42] = 32'b00000001010000100001000110000011; // 0x01421183 | lh   x3, 20(x4)
      Imemory[43] = 32'b00000000000000101001011000000011; // 0x00029503 | lh   x6, 0(x5)
      Imemory[44] = 32'b00000110010000100100000110000011; // 0x06422183 | lw   x3, 100(x4)
      Imemory[45] = 32'b11111111100000101010011000000011; // 0xff82b603 | lw   x6, -8(x5)
      Imemory[46] = 32'b00000001100100000000100110000011; // 0x01900183 | lbu  x3, 25(x1)
      Imemory[47] = 32'b11111111111000010000111000000011; // 0xffe10703 | lbu  x6, -2(x2)
      Imemory[48] = 32'b00000011001000100101100110000011; // 0x03229583 | lhu  x3, 50(x4)
      Imemory[49] = 32'b00000000010000000001111000000011; // 0x00400783 | lhu  x6, 4(x1)

      // ===== JALR đảm bảo PC tuần tự +4: auipc x1,0; addi x1,x1,4; jalr x3,x1,0 =====
      Imemory[50] = 32'b00000000000000000000_00001_0010111;     // 0x00000097 | auipc x1, 0        | x1 = PC
		Imemory[51] = 32'b00000000100000001000000111100111;   // 0x00c081e7 | jalr  x3, x1, 8   | PC = (x1 + 8) & ~1 = PC + 4
		Imemory[52] = 32'b000000000000_00000_000_00000_0010011;   // 0x00000013 | addi  x0, x0, 0    | nop giữ chỗ (đảm bảo tổng 76 lệnh)

      // ===== S-type (giống R-type: rs1, rs2 ∈ {x1,x2,x4,x5}) =====
      Imemory[53] = 32'b00000000000100010000011110100011; // 0x001107a3 | sb   x1, 15(x2)
      Imemory[54] = 32'b11111110011100100000111010100011; // 0xfe720ea3 | sb   x5, -3(x4)
      Imemory[55] = 32'b00000000001100010001111100100011; // 0x00311f23 | sh   x1, 30(x2)
      Imemory[56] = 32'b00000000010100100001000000100011; // 0x00521023 | sh   x5, 0(x4)
      Imemory[57] = 32'b00001100001000101010010000100011; // 0x00a2c223 | sw   x2, 200(x5)
      Imemory[58] = 32'b11111110010000010010101000100011; // 0xfec14a23 | sw   x4, -12(x2)

      // ===== B-type (tất cả imm = 4) =====
      Imemory[59] = 32'b00000000001000001000001001100011; // 0x00208263 | beq  x1,  x2, 4
      Imemory[60] = 32'b00000001001101000100001001100011; // 0x01344263 | beq  x8,  x9, 4
      Imemory[61] = 32'b00000000010000011001001001100011; // 0x00419263 | bne  x3,  x4, 4
      Imemory[62] = 32'b00000001010101010001001001100011; // 0x01554263 | bne  x10, x11, 4
      Imemory[63] = 32'b00000000011000101100001001100011; // 0x0062c263 | blt  x5,  x6, 4
      Imemory[64] = 32'b00000001110101100100001001100011; // 0x01d64263 | blt  x12, x13, 4
      Imemory[65] = 32'b00000000100000111101001001100011; // 0x0083d263 | bge  x7,  x8, 4
      Imemory[66] = 32'b00000001111001111101001001100011; // 0x01e7d263 | bge  x14, x15, 4
      Imemory[67] = 32'b00000000001100001110001001100011; // 0x0030e263 | bltu x1,  x3, 4
      Imemory[68] = 32'b00000001001001001110001001100011; // 0x0124e263 | bltu x9,  x10, 4
      Imemory[69] = 32'b00000000101000100111001001100011; // 0x00a27763 | bgeu x4,  x5, 4
      Imemory[70] = 32'b00000001100001100111001001100011; // 0x01867763 | bgeu x11, x12, 4

      // ===== U-type (giữ nguyên) =====
      Imemory[71] = 32'b00010010001101000101000010110111; // 0x123450b7 | lui   x1, 0x12345
      Imemory[72] = 32'b10101011110011011110010000110111; // 0xabcde437 | lui   x8, 0xABCDE
      Imemory[73] = 32'b00000001000000000000000100010111; // 0x01000117 | auipc x2, 0x1000
		Imemory[74] = 32'b00000101011001111000010010010111; // 0x05678497 | auipc x9, 0x5678
		

      // ===== J-type (imm = 4 để PC tiến +4) =====
      Imemory[75] = 32'b00000000000000000001000011101111; // 0x004001ef | jal   x3, 4
		
      
      
    end
  end
  
endmodule