    initial begin
        // Expected results for 51 instructions that write to registers

        expected_pcs[ 0]  = 0x00000004; expected_results[ 0]  = 32'h00000030; expected_rds[ 0]  = 5'd 3;
        expected_pcs[ 1]  = 0x00000008; expected_results[ 1]  = 32'hfffffff0; expected_rds[ 1]  = 5'd12;
        expected_pcs[ 2]  = 0x0000000c; expected_results[ 2]  = 32'h00000010; expected_rds[ 2]  = 5'd 3;
        expected_pcs[ 3]  = 0x00000010; expected_results[ 3]  = 32'h00000001; expected_rds[ 3]  = 5'd12;
        expected_pcs[ 4]  = 0x00000014; expected_results[ 4]  = 32'h00000000; expected_rds[ 4]  = 5'd 3;
        expected_pcs[ 5]  = 0x00000018; expected_results[ 5]  = 32'h00000040; expected_rds[ 5]  = 5'd12;
        expected_pcs[ 6]  = 0x0000001c; expected_results[ 6]  = 32'h00000040; expected_rds[ 6]  = 5'd 3;
        expected_pcs[ 7]  = 0x00000020; expected_results[ 7]  = 32'h00000000; expected_rds[ 7]  = 5'd12;
        expected_pcs[ 8]  = 0x00000024; expected_results[ 8]  = 32'h00000050; expected_rds[ 8]  = 5'd 3;
        expected_pcs[ 9]  = 0x00000028; expected_results[ 9]  = 32'h00000000; expected_rds[ 9]  = 5'd12;
        expected_pcs[10]  = 0x0000002c; expected_results[10]  = 32'h00000010; expected_rds[10]  = 5'd12;
        expected_pcs[11]  = 0x00000030; expected_results[11]  = 32'h00000010; expected_rds[11]  = 5'd 3;
        expected_pcs[12]  = 0x00000034; expected_results[12]  = 32'h00000020; expected_rds[12]  = 5'd12;
        expected_pcs[13]  = 0x00000038; expected_results[13]  = 32'h00000001; expected_rds[13]  = 5'd 3;
        expected_pcs[14]  = 0x0000003c; expected_results[14]  = 32'h00000050; expected_rds[14]  = 5'd12;
        expected_pcs[15]  = 0x00000040; expected_results[15]  = 32'h00000060; expected_rds[15]  = 5'd 3;
        expected_pcs[16]  = 0x00000044; expected_results[16]  = 32'h00000000; expected_rds[16]  = 5'd12;
        expected_pcs[17]  = 0x00000048; expected_results[17]  = 32'h00000050; expected_rds[17]  = 5'd 3;
        expected_pcs[18]  = 0x0000004c; expected_results[18]  = 32'h00000060; expected_rds[18]  = 5'd12;
        expected_pcs[19]  = 0x00000050; expected_results[19]  = 32'h00000010; expected_rds[19]  = 5'd 3;
        expected_pcs[20]  = 0x00000054; expected_results[20]  = 32'h0000001c; expected_rds[20]  = 5'd 3;
        expected_pcs[21]  = 0x00000058; expected_results[21]  = 32'hffffffee; expected_rds[21]  = 5'd12;
        expected_pcs[22]  = 0x0000005c; expected_results[22]  = 32'h00000000; expected_rds[22]  = 5'd 3;
        expected_pcs[23]  = 0x00000060; expected_results[23]  = 32'h00000000; expected_rds[23]  = 5'd12;
        expected_pcs[24]  = 0x00000064; expected_results[24]  = 32'h00000001; expected_rds[24]  = 5'd12;
        expected_pcs[25]  = 0x00000068; expected_results[25]  = 32'h00000000; expected_rds[25]  = 5'd 3;
        expected_pcs[26]  = 0x0000006c; expected_results[26]  = 32'h0000005f; expected_rds[26]  = 5'd12;
        expected_pcs[27]  = 0x00000070; expected_results[27]  = 32'h00000045; expected_rds[27]  = 5'd 3;
        expected_pcs[28]  = 0x00000074; expected_results[28]  = 32'h00000010; expected_rds[28]  = 5'd 3;
        expected_pcs[29]  = 0x00000078; expected_results[29]  = 32'h00000028; expected_rds[29]  = 5'd12;
        expected_pcs[30]  = 0x0000007c; expected_results[30]  = 32'h00000000; expected_rds[30]  = 5'd12;
        expected_pcs[31]  = 0x00000080; expected_results[31]  = 32'h00000000; expected_rds[31]  = 5'd19;
        expected_pcs[32]  = 0x00000084; expected_results[32]  = 32'h00000080; expected_rds[32]  = 5'd 3;
        expected_pcs[33]  = 0x00000088; expected_results[33]  = 32'h00002000; expected_rds[33]  = 5'd12;
        expected_pcs[34]  = 0x0000008c; expected_results[34]  = 32'h00000005; expected_rds[34]  = 5'd 3;
        expected_pcs[35]  = 0x00000090; expected_results[35]  = 32'h00000000; expected_rds[35]  = 5'd12;
        expected_pcs[36]  = 0x00000094; expected_results[36]  = 32'h00000010; expected_rds[36]  = 5'd 3;
        expected_pcs[37]  = 0x00000098; expected_results[37]  = 32'h00000000; expected_rds[37]  = 5'd12;
        expected_pcs[38]  = 0x0000009c; expected_results[38]  = 32'h00000050; expected_rds[38]  = 5'd 3;
        expected_pcs[39]  = 0x000000a0; expected_results[39]  = 32'h00000000; expected_rds[39]  = 5'd 3;
        expected_pcs[40]  = 0x000000a8; expected_results[40]  = 32'h00000000; expected_rds[40]  = 5'd 3;
        expected_pcs[41]  = 0x000000ac; expected_results[41]  = 32'h00000000; expected_rds[41]  = 5'd12;
        expected_pcs[42]  = 0x000000b0; expected_results[42]  = 32'h00000000; expected_rds[42]  = 5'd 3;
        expected_pcs[43]  = 0x000000b4; expected_results[43]  = 32'h00000000; expected_rds[43]  = 5'd12;
        expected_pcs[44]  = 0x000000b8; expected_results[44]  = 32'h00000000; expected_rds[44]  = 5'd19;
        expected_pcs[45]  = 0x000000bc; expected_results[45]  = 32'h00000000; expected_rds[45]  = 5'd28;
        expected_pcs[46]  = 0x000000c0; expected_results[46]  = 32'h00000000; expected_rds[46]  = 5'd19;
        expected_pcs[47]  = 0x00000114; expected_results[47]  = 32'habcde000; expected_rds[47]  = 5'd 8;
        expected_pcs[48]  = 0x00000118; expected_results[48]  = 32'h01000118; expected_rds[48]  = 5'd 2;
        expected_pcs[49]  = 0x0000011c; expected_results[49]  = 32'h0567811c; expected_rds[49]  = 5'd 9;
        expected_pcs[50]  = 0x00000120; expected_results[50]  = 32'h00000124; expected_rds[50]  = 5'd 1;
    end