// =============================================================================
// Sequence: TC 6.2.2 - STORE_HALF_MASK Instruction
// =============================================================================
// Category: Memory System
// Priority: HIGH
// Description: SH halfword masking
// =============================================================================

class tc_6_2_2_store_half_mask_seq extends uvm_sequence #(rv32i_transaction);
    
    `uvm_object_utils(tc_6_2_2_store_half_mask_seq)
    
    function new(string name = "tc_6_2_2_store_half_mask_seq");
        super.new(name);
    endfunction
    
    task body();
        rv32i_transaction tr;
        
        `uvm_info(get_type_name(), "Starting STORE_HALF_MASK sequence", UVM_MEDIUM)
        
        // ======================================================================
        // Test Case: STORE_HALF_MASK - SH halfword masking
        // ======================================================================
        tr = rv32i_transaction::type_id::create("store_half_mask_test");
        start_item(tr);
        
        tr.test_name = "STORE_HALF_MASK Test";
        // TODO: Configure instruction encoding and test values
        // tr.opcode = ...;
        // tr.funct3 = ...;
        // tr.rd = ...;
        // tr.rs1 = ...;
        // tr.rs2 = ...;
        // tr.instruction = {tr.funct7, tr.rs2, tr.rs1, tr.funct3, tr.rd, tr.opcode};
        
        finish_item(tr);
        `uvm_info(get_type_name(), "Sent: STORE_HALF_MASK test transaction", UVM_HIGH)
        
        `uvm_info(get_type_name(), "STORE_HALF_MASK sequence completed", UVM_MEDIUM)
        
    endtask

endclass : tc_6_2_2_store_half_mask_seq
