// =============================================================================
// Test Package
// =============================================================================
// Contains all test classes organized by priority
// =============================================================================

package test_pkg;

    import uvm_pkg::*;
    import component_pkg::*;
    import seq_pkg::*;
    `include "uvm_macros.svh"

    // Base test
    `include "tests/base_test.sv"

    // ==========================================================================
    // Golden Verification Tests (37 tests)
    // ==========================================================================
    `include "tests/golden_verification/tc_1_1_10_and_golden_test.sv"
    `include "tests/golden_verification/tc_1_1_1_add_golden_test.sv"
    `include "tests/golden_verification/tc_1_1_2_sub_golden_test.sv"
    `include "tests/golden_verification/tc_1_1_3_sll_golden_test.sv"
    `include "tests/golden_verification/tc_1_1_4_slt_golden_test.sv"
    `include "tests/golden_verification/tc_1_1_5_sltu_golden_test.sv"
    `include "tests/golden_verification/tc_1_1_6_xor_golden_test.sv"
    `include "tests/golden_verification/tc_1_1_7_srl_golden_test.sv"
    `include "tests/golden_verification/tc_1_1_8_sra_golden_test.sv"
    `include "tests/golden_verification/tc_1_1_9_or_golden_test.sv"
    `include "tests/golden_verification/tc_1_2_1_addi_golden_test.sv"
    `include "tests/golden_verification/tc_1_2_2_slti_golden_test.sv"
    `include "tests/golden_verification/tc_1_2_3_sltiu_golden_test.sv"
    `include "tests/golden_verification/tc_1_2_4_xori_golden_test.sv"
    `include "tests/golden_verification/tc_1_2_5_ori_golden_test.sv"
    `include "tests/golden_verification/tc_1_2_6_andi_golden_test.sv"
    `include "tests/golden_verification/tc_1_2_7_slli_golden_test.sv"
    `include "tests/golden_verification/tc_1_2_8_srli_golden_test.sv"
    `include "tests/golden_verification/tc_1_2_9_srai_golden_test.sv"
    `include "tests/golden_verification/tc_1_3_1_lw_golden_test.sv"
    `include "tests/golden_verification/tc_1_3_2_lh_golden_test.sv"
    `include "tests/golden_verification/tc_1_3_3_lhu_golden_test.sv"
    `include "tests/golden_verification/tc_1_3_4_lb_golden_test.sv"
    `include "tests/golden_verification/tc_1_3_5_lbu_golden_test.sv"
    `include "tests/golden_verification/tc_1_4_1_sw_golden_test.sv"
    `include "tests/golden_verification/tc_1_4_2_sh_golden_test.sv"
    `include "tests/golden_verification/tc_1_4_3_sb_golden_test.sv"
    `include "tests/golden_verification/tc_1_5_1_beq_golden_test.sv"
    `include "tests/golden_verification/tc_1_5_2_bne_golden_test.sv"
    `include "tests/golden_verification/tc_1_5_3_blt_golden_test.sv"
    `include "tests/golden_verification/tc_1_5_4_bge_golden_test.sv"
    `include "tests/golden_verification/tc_1_5_5_bltu_golden_test.sv"
    `include "tests/golden_verification/tc_1_5_6_bgeu_golden_test.sv"
    `include "tests/golden_verification/tc_1_6_1_jal_golden_test.sv"
    `include "tests/golden_verification/tc_1_6_2_jalr_golden_test.sv"
    `include "tests/golden_verification/tc_1_7_1_lui_golden_test.sv"
    `include "tests/golden_verification/tc_1_7_2_auipc_golden_test.sv"

    // ==========================================================================
    // Critical Priority Tests (78 tests)
    // ==========================================================================
    `include "tests/critical/tc_1_1_10_and_test.sv"
    `include "tests/critical/tc_1_1_1_add_test.sv"
    `include "tests/critical/tc_1_1_2_sub_test.sv"
    `include "tests/critical/tc_1_1_3_sll_test.sv"
    `include "tests/critical/tc_1_1_4_slt_test.sv"
    `include "tests/critical/tc_1_1_5_sltu_test.sv"
    `include "tests/critical/tc_1_1_6_xor_test.sv"
    `include "tests/critical/tc_1_1_7_srl_test.sv"
    `include "tests/critical/tc_1_1_8_sra_test.sv"
    `include "tests/critical/tc_1_1_9_or_test.sv"
    `include "tests/critical/tc_1_2_1_addi_test.sv"
    `include "tests/critical/tc_1_2_2_slti_test.sv"
    `include "tests/critical/tc_1_2_3_sltiu_test.sv"
    `include "tests/critical/tc_1_2_4_xori_test.sv"
    `include "tests/critical/tc_1_2_5_ori_test.sv"
    `include "tests/critical/tc_1_2_6_andi_test.sv"
    `include "tests/critical/tc_1_2_7_slli_test.sv"
    `include "tests/critical/tc_1_2_8_srli_test.sv"
    `include "tests/critical/tc_1_2_9_srai_test.sv"
    `include "tests/critical/tc_1_3_1_lw_test.sv"
    `include "tests/critical/tc_1_3_2_lh_test.sv"
    `include "tests/critical/tc_1_3_3_lhu_test.sv"
    `include "tests/critical/tc_1_3_4_lb_test.sv"
    `include "tests/critical/tc_1_3_5_lbu_test.sv"
    `include "tests/critical/tc_1_4_1_sw_test.sv"
    `include "tests/critical/tc_1_4_2_sh_test.sv"
    `include "tests/critical/tc_1_4_3_sb_test.sv"
    `include "tests/critical/tc_1_5_1_beq_test.sv"
    `include "tests/critical/tc_1_5_2_bne_test.sv"
    `include "tests/critical/tc_1_5_3_blt_test.sv"
    `include "tests/critical/tc_1_5_4_bge_test.sv"
    `include "tests/critical/tc_1_5_5_bltu_test.sv"
    `include "tests/critical/tc_1_5_6_bgeu_test.sv"
    `include "tests/critical/tc_1_6_1_jal_test.sv"
    `include "tests/critical/tc_1_6_2_jalr_test.sv"
    `include "tests/critical/tc_1_7_1_lui_test.sv"
    `include "tests/critical/tc_1_7_2_auipc_test.sv"
    `include "tests/critical/tc_2_1_1_raw_ex_ex_test.sv"
    `include "tests/critical/tc_2_1_2_raw_mem_ex_test.sv"
    `include "tests/critical/tc_2_1_3_raw_wb_ex_test.sv"
    `include "tests/critical/tc_2_1_4_raw_double_test.sv"
    `include "tests/critical/tc_2_2_1_load_use_stall_test.sv"
    `include "tests/critical/tc_2_2_2_load_forward_test.sv"
    `include "tests/critical/tc_2_2_3_back_to_back_loads_test.sv"
    `include "tests/critical/tc_2_3_1_rs1_forward_test.sv"
    `include "tests/critical/tc_2_3_2_rs2_forward_test.sv"
    `include "tests/critical/tc_2_3_3_both_rs_forward_test.sv"
    `include "tests/critical/tc_2_3_4_store_data_forward_test.sv"
    `include "tests/critical/tc_2_4_1_chain_raw_test.sv"
    `include "tests/critical/tc_2_4_2_multiple_consumers_test.sv"
    `include "tests/critical/tc_2_4_3_interleaved_hazards_test.sv"
    `include "tests/critical/tc_2_5_1_x0_raw_test.sv"
    `include "tests/critical/tc_2_5_2_x0_write_ignored_test.sv"
    `include "tests/critical/tc_3_1_1_branch_taken_test.sv"
    `include "tests/critical/tc_3_1_2_branch_not_taken_test.sv"
    `include "tests/critical/tc_3_1_3_backward_branch_test.sv"
    `include "tests/critical/tc_3_1_4_forward_branch_test.sv"
    `include "tests/critical/tc_3_2_1_jal_forward_test.sv"
    `include "tests/critical/tc_3_2_2_jal_backward_test.sv"
    `include "tests/critical/tc_3_2_3_jalr_computed_test.sv"
    `include "tests/critical/tc_3_2_4_jalr_return_test.sv"
    `include "tests/critical/tc_3_3_1_branch_after_load_test.sv"
    `include "tests/critical/tc_3_3_2_branch_with_forward_test.sv"
    `include "tests/critical/tc_3_3_3_jump_after_alu_test.sv"
    `include "tests/critical/tc_3_4_1_back_to_back_branches_test.sv"
    `include "tests/critical/tc_3_4_2_nested_branches_test.sv"
    `include "tests/critical/tc_3_4_3_branch_in_delay_test.sv"
    `include "tests/critical/tc_3_5_1_flush_if_test.sv"
    `include "tests/critical/tc_3_5_2_flush_id_test.sv"
    `include "tests/critical/tc_9_1_1_ex_to_ex_rs1_test.sv"
    `include "tests/critical/tc_9_1_2_ex_to_ex_rs2_test.sv"
    `include "tests/critical/tc_9_1_3_ex_to_ex_both_test.sv"
    `include "tests/critical/tc_9_2_1_mem_to_ex_rs1_test.sv"
    `include "tests/critical/tc_9_2_2_mem_to_ex_rs2_test.sv"
    `include "tests/critical/tc_9_2_3_mem_to_ex_both_test.sv"
    `include "tests/critical/tc_9_3_1_load_forward_test.sv"
    `include "tests/critical/tc_9_3_2_alu_to_branch_test.sv"
    `include "tests/critical/tc_9_3_3_alu_to_store_test.sv"

    // ==========================================================================
    // High Priority Tests (50 tests)
    // ==========================================================================
    `include "tests/high/tc_12_1_1_jal_return_addr_test.sv"
    `include "tests/high/tc_12_1_2_jalr_return_addr_test.sv"
    `include "tests/high/tc_12_2_1_jal_to_x0_test.sv"
    `include "tests/high/tc_12_2_2_jalr_to_x0_test.sv"
    `include "tests/high/tc_4_1_1_overflow_add_test.sv"
    `include "tests/high/tc_4_1_2_underflow_sub_test.sv"
    `include "tests/high/tc_4_1_3_max_shift_test.sv"
    `include "tests/high/tc_4_2_1_x0_read_test.sv"
    `include "tests/high/tc_4_2_2_x0_write_test.sv"
    `include "tests/high/tc_4_2_3_x0_both_test.sv"
    `include "tests/high/tc_4_3_1_max_pos_imm_test.sv"
    `include "tests/high/tc_4_3_2_max_neg_imm_test.sv"
    `include "tests/high/tc_4_3_3_zero_imm_test.sv"
    `include "tests/high/tc_4_4_1_mem_addr_0_test.sv"
    `include "tests/high/tc_4_4_2_mem_addr_max_test.sv"
    `include "tests/high/tc_4_4_3_mem_unaligned_test.sv"
    `include "tests/high/tc_4_5_1_branch_target_0_test.sv"
    `include "tests/high/tc_4_5_2_branch_self_test.sv"
    `include "tests/high/tc_4_5_3_branch_max_offset_test.sv"
    `include "tests/high/tc_4_6_1_all_ones_test.sv"
    `include "tests/high/tc_4_6_2_all_zeros_test.sv"
    `include "tests/high/tc_4_6_3_alternating_bits_test.sv"
    `include "tests/high/tc_4_6_4_single_bit_test.sv"
    `include "tests/high/tc_5_1_1_raw_and_branch_test.sv"
    `include "tests/high/tc_5_1_2_load_use_and_branch_test.sv"
    `include "tests/high/tc_5_1_3_forward_and_jump_test.sv"
    `include "tests/high/tc_5_2_1_loop_with_hazards_test.sv"
    `include "tests/high/tc_5_2_2_nested_loops_test.sv"
    `include "tests/high/tc_5_2_3_loop_unroll_test.sv"
    `include "tests/high/tc_5_3_1_function_call_test.sv"
    `include "tests/high/tc_5_3_2_function_return_test.sv"
    `include "tests/high/tc_5_3_3_nested_calls_test.sv"
    `include "tests/high/tc_5_4_1_mixed_hazards_test.sv"
    `include "tests/high/tc_6_1_1_load_byte_sign_ext_test.sv"
    `include "tests/high/tc_6_1_2_load_byte_zero_ext_test.sv"
    `include "tests/high/tc_6_1_3_load_half_sign_ext_test.sv"
    `include "tests/high/tc_6_1_4_load_half_zero_ext_test.sv"
    `include "tests/high/tc_6_2_1_store_byte_mask_test.sv"
    `include "tests/high/tc_6_2_2_store_half_mask_test.sv"
    `include "tests/high/tc_6_2_3_store_word_test.sv"
    `include "tests/high/tc_6_3_1_load_word_align_test.sv"
    `include "tests/high/tc_6_3_2_load_half_align_test.sv"
    `include "tests/high/tc_6_3_3_store_align_test.sv"
    `include "tests/high/tc_6_4_1_load_store_same_addr_test.sv"
    `include "tests/high/tc_6_4_2_store_load_forward_test.sv"
    `include "tests/high/tc_6_4_3_back_to_back_mem_test.sv"
    `include "tests/high/tc_6_5_1_mem_offset_pos_test.sv"
    `include "tests/high/tc_6_5_2_mem_offset_neg_test.sv"
    `include "tests/high/tc_6_5_3_mem_offset_zero_test.sv"
    `include "tests/high/tc_6_5_4_mem_offset_max_test.sv"

    // ==========================================================================
    // Medium Priority Tests (27 tests)
    // ==========================================================================
    `include "tests/medium/tc_11_1_1_add_overflow_pos_test.sv"
    `include "tests/medium/tc_11_1_2_add_overflow_neg_test.sv"
    `include "tests/medium/tc_11_1_3_sub_underflow_test.sv"
    `include "tests/medium/tc_11_2_1_slt_edge_cases_test.sv"
    `include "tests/medium/tc_11_2_2_sltu_edge_cases_test.sv"
    `include "tests/medium/tc_11_2_3_shift_edge_cases_test.sv"
    `include "tests/medium/tc_13_1_1_imm_12bit_max_test.sv"
    `include "tests/medium/tc_13_1_2_imm_20bit_max_test.sv"
    `include "tests/medium/tc_13_1_3_imm_sign_ext_test.sv"
    `include "tests/medium/tc_13_1_4_imm_zero_ext_test.sv"
    `include "tests/medium/tc_14_1_1_long_sequence_test.sv"
    `include "tests/medium/tc_14_1_2_deep_nesting_test.sv"
    `include "tests/medium/tc_14_1_3_max_dependencies_test.sv"
    `include "tests/medium/tc_7_1_1_all_regs_write_test.sv"
    `include "tests/medium/tc_7_1_2_all_regs_read_test.sv"
    `include "tests/medium/tc_7_2_1_x0_always_zero_test.sv"
    `include "tests/medium/tc_7_2_2_x0_as_source_test.sv"
    `include "tests/medium/tc_7_3_1_same_reg_src_dst_test.sv"
    `include "tests/medium/tc_7_3_2_all_same_reg_test.sv"
    `include "tests/medium/tc_7_4_1_rapid_reuse_test.sv"
    `include "tests/medium/tc_7_4_2_reg_ping_pong_test.sv"
    `include "tests/medium/tc_8_1_1_single_stall_test.sv"
    `include "tests/medium/tc_8_1_2_multi_stall_test.sv"
    `include "tests/medium/tc_8_2_1_stall_recovery_test.sv"
    `include "tests/medium/tc_8_2_2_stall_then_branch_test.sv"
    `include "tests/medium/tc_8_3_1_back_to_back_stalls_test.sv"
    `include "tests/medium/tc_8_3_2_stall_patterns_test.sv"

    // ==========================================================================
    // Low Priority Tests (3 tests)
    // ==========================================================================
    `include "tests/low/tc_10_1_1_cpi_no_hazards_test.sv"
    `include "tests/low/tc_10_1_2_cpi_with_hazards_test.sv"
    `include "tests/low/tc_10_1_3_cpi_worst_case_test.sv"

endpackage : test_pkg
