// =============================================================================
// Sequence: TC 3.3.3 - JUMP_AFTER_ALU Instruction
// =============================================================================
// Category: Control Hazards
// Priority: CRITICAL
// Description: Jump after ALU operation
// =============================================================================

class tc_3_3_3_jump_after_alu_seq extends uvm_sequence #(rv32i_transaction);
    
    `uvm_object_utils(tc_3_3_3_jump_after_alu_seq)
    
    function new(string name = "tc_3_3_3_jump_after_alu_seq");
        super.new(name);
    endfunction
    
    task body();
        rv32i_transaction tr;
        
        `uvm_info(get_type_name(), "Starting JUMP_AFTER_ALU sequence", UVM_MEDIUM)
        
        // ======================================================================
        // Test Case: JUMP_AFTER_ALU - Jump after ALU operation
        // ======================================================================
        tr = rv32i_transaction::type_id::create("jump_after_alu_test");
        start_item(tr);
        
        tr.test_name = "JUMP_AFTER_ALU Test";
        // TODO: Configure instruction encoding and test values
        // tr.opcode = ...;
        // tr.funct3 = ...;
        // tr.rd = ...;
        // tr.rs1 = ...;
        // tr.rs2 = ...;
        // tr.instruction = {tr.funct7, tr.rs2, tr.rs1, tr.funct3, tr.rd, tr.opcode};
        
        finish_item(tr);
        `uvm_info(get_type_name(), "Sent: JUMP_AFTER_ALU test transaction", UVM_HIGH)
        
        `uvm_info(get_type_name(), "JUMP_AFTER_ALU sequence completed", UVM_MEDIUM)
        
    endtask

endclass : tc_3_3_3_jump_after_alu_seq
