// =============================================================================
// Sequence: TC 1.7.1 - LUI Instruction
// =============================================================================
// Category: ISA Coverage
// Priority: CRITICAL
// Description: Load upper immediate
// =============================================================================

class tc_1_7_1_lui_seq extends uvm_sequence #(rv32i_transaction);
    
    `uvm_object_utils(tc_1_7_1_lui_seq)
    
    function new(string name = "tc_1_7_1_lui_seq");
        super.new(name);
    endfunction
    
    task body();
        rv32i_transaction tr;
        
        `uvm_info(get_type_name(), "Starting LUI sequence", UVM_MEDIUM)
        
        // ======================================================================
        // Test Case: LUI - Load upper immediate
        // ======================================================================
        tr = rv32i_transaction::type_id::create("lui_test");
        start_item(tr);
        
        tr.test_name = "LUI Test";
        // TODO: Configure instruction encoding and test values
        // tr.opcode = ...;
        // tr.funct3 = ...;
        // tr.rd = ...;
        // tr.rs1 = ...;
        // tr.rs2 = ...;
        // tr.instruction = {tr.funct7, tr.rs2, tr.rs1, tr.funct3, tr.rd, tr.opcode};
        
        finish_item(tr);
        `uvm_info(get_type_name(), "Sent: LUI test transaction", UVM_HIGH)
        
        `uvm_info(get_type_name(), "LUI sequence completed", UVM_MEDIUM)
        
    endtask

endclass : tc_1_7_1_lui_seq
