// =============================================================================
// Test Case 8.3.2: STALL_PATTERNS
// =============================================================================
// Category: Pipeline Stalls
// Priority: MEDIUM
// Description: Various stall patterns
// =============================================================================

class tc_8_3_2_stall_patterns_test extends base_test;
    
    `uvm_component_utils(tc_8_3_2_stall_patterns_test)
    
    function new(string name = "tc_8_3_2_stall_patterns_test", uvm_component parent = null);
        super.new(name, parent);
    endfunction
    
    function void build_phase(uvm_phase phase);
        super.build_phase(phase);
        
        // Override golden log file for this test
        golden_log_file = "tests/golden/tc_8_3_2_stall_patterns_golden.log";
        uvm_config_db#(string)::set(this, "env.scoreboard.golden", 
                                    "golden_log_file", golden_log_file);
    endfunction
    
    task run_phase(uvm_phase phase);
        tc_8_3_2_stall_patterns_seq seq;
        
        phase.raise_objection(this);
        
        `uvm_info(get_type_name(), "\n=== Starting TC 8.3.2: STALL_PATTERNS ===", UVM_LOW)
        
        // Create and start sequence
        seq = tc_8_3_2_stall_patterns_seq::type_id::create("seq");
        seq.start(env.agent.sequencer);
        
        // Wait for completion
        #1000;
        
        `uvm_info(get_type_name(), "=== TC 8.3.2: STALL_PATTERNS Complete ===\n", UVM_LOW)
        
        phase.drop_objection(this);
    endtask

endclass : tc_8_3_2_stall_patterns_test
