// =============================================================================
// Sequence: TC 1.1.5 - SLTU Instruction
// =============================================================================
// Category: ISA Coverage
// Priority: CRITICAL
// Description: Set less than (unsigned)
// =============================================================================

class tc_1_1_5_sltu_seq extends uvm_sequence #(rv32i_transaction);
    
    `uvm_object_utils(tc_1_1_5_sltu_seq)
    
    function new(string name = "tc_1_1_5_sltu_seq");
        super.new(name);
    endfunction
    
    task body();
        rv32i_transaction tr;
        
        `uvm_info(get_type_name(), "Starting SLTU sequence", UVM_MEDIUM)
        
        // ======================================================================
        // Test Case: SLTU - Set less than (unsigned)
        // ======================================================================
        tr = rv32i_transaction::type_id::create("sltu_test");
        start_item(tr);
        
        tr.test_name = "SLTU Test";
        // TODO: Configure instruction encoding and test values
        // tr.opcode = ...;
        // tr.funct3 = ...;
        // tr.rd = ...;
        // tr.rs1 = ...;
        // tr.rs2 = ...;
        // tr.instruction = {tr.funct7, tr.rs2, tr.rs1, tr.funct3, tr.rd, tr.opcode};
        
        finish_item(tr);
        `uvm_info(get_type_name(), "Sent: SLTU test transaction", UVM_HIGH)
        
        `uvm_info(get_type_name(), "SLTU sequence completed", UVM_MEDIUM)
        
    endtask

endclass : tc_1_1_5_sltu_seq
