// =============================================================================
// Sequence: TC 1.1.2 - SUB Instruction
// =============================================================================
// Category: ISA Coverage
// Priority: CRITICAL
// Description: Basic subtraction
// =============================================================================

class tc_1_1_2_sub_seq extends uvm_sequence #(rv32i_transaction);
    
    `uvm_object_utils(tc_1_1_2_sub_seq)
    
    function new(string name = "tc_1_1_2_sub_seq");
        super.new(name);
    endfunction
    
    task body();
        rv32i_transaction tr;
        
        `uvm_info(get_type_name(), "Starting SUB sequence", UVM_MEDIUM)
        
        // ======================================================================
        // Test Case: SUB - Basic subtraction
        // ======================================================================
        tr = rv32i_transaction::type_id::create("sub_test");
        start_item(tr);
        
        tr.test_name = "SUB Test";
        // TODO: Configure instruction encoding and test values
        // tr.opcode = ...;
        // tr.funct3 = ...;
        // tr.rd = ...;
        // tr.rs1 = ...;
        // tr.rs2 = ...;
        // tr.instruction = {tr.funct7, tr.rs2, tr.rs1, tr.funct3, tr.rd, tr.opcode};
        
        finish_item(tr);
        `uvm_info(get_type_name(), "Sent: SUB test transaction", UVM_HIGH)
        
        `uvm_info(get_type_name(), "SUB sequence completed", UVM_MEDIUM)
        
    endtask

endclass : tc_1_1_2_sub_seq
