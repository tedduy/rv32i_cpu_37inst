// =============================================================================
// Test Case 15.1.3: MAX_DEPENDENCIES
// =============================================================================
// Category: Stress Tests
// Priority: MEDIUM
// Description: Maximum dependency chains
// =============================================================================

class tc_15_1_3_max_dependencies_test extends base_test;
    
    `uvm_component_utils(tc_15_1_3_max_dependencies_test)
    
    function new(string name = "tc_15_1_3_max_dependencies_test", uvm_component parent = null);
        super.new(name, parent);
    endfunction
    
    function void build_phase(uvm_phase phase);
        super.build_phase(phase);
        
        // Override spike log file for this test
        spike_log_file = "tests/golden/tc_15_1_3_max_dependencies_spike.log";
        uvm_config_db#(string)::set(this, "env.scoreboard.spike", 
                                    "spike_log_file", spike_log_file);
    endfunction
    
    task run_phase(uvm_phase phase);
        tc_15_1_3_max_dependencies_seq seq;
        
        phase.raise_objection(this);
        
        `uvm_info(get_type_name(), "\n=== Starting TC 15.1.3: MAX_DEPENDENCIES ===", UVM_LOW)
        
        // Create and start sequence
        seq = tc_15_1_3_max_dependencies_seq::type_id::create("seq");
        seq.start(env.agent.sequencer);
        
        // Wait for completion
        #1000;
        
        `uvm_info(get_type_name(), "=== TC 15.1.3: MAX_DEPENDENCIES Complete ===\n", UVM_LOW)
        
        phase.drop_objection(this);
    endtask

endclass : tc_15_1_3_max_dependencies_test
