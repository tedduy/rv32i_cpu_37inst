// =============================================================================
// Sequence: TC 2.4.1 - CHAIN_RAW Instruction
// =============================================================================
// Category: Data Hazards
// Priority: CRITICAL
// Description: Chain of RAW dependencies
// =============================================================================

class tc_2_4_1_chain_raw_seq extends uvm_sequence #(rv32i_transaction);
    
    `uvm_object_utils(tc_2_4_1_chain_raw_seq)
    
    function new(string name = "tc_2_4_1_chain_raw_seq");
        super.new(name);
    endfunction
    
    task body();
        rv32i_transaction tr;
        
        `uvm_info(get_type_name(), "Starting CHAIN_RAW sequence", UVM_MEDIUM)
        
        // ======================================================================
        // Test Case: CHAIN_RAW - Chain of RAW dependencies
        // ======================================================================
        tr = rv32i_transaction::type_id::create("chain_raw_test");
        start_item(tr);
        
        tr.test_name = "CHAIN_RAW Test";
        // TODO: Configure instruction encoding and test values
        // tr.opcode = ...;
        // tr.funct3 = ...;
        // tr.rd = ...;
        // tr.rs1 = ...;
        // tr.rs2 = ...;
        // tr.instruction = {tr.funct7, tr.rs2, tr.rs1, tr.funct3, tr.rd, tr.opcode};
        
        finish_item(tr);
        `uvm_info(get_type_name(), "Sent: CHAIN_RAW test transaction", UVM_HIGH)
        
        `uvm_info(get_type_name(), "CHAIN_RAW sequence completed", UVM_MEDIUM)
        
    endtask

endclass : tc_2_4_1_chain_raw_seq
