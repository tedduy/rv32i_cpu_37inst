// =============================================================================
// Sequence: TC 1.1.8 - SRA Instruction
// =============================================================================
// Category: ISA Coverage
// Priority: CRITICAL
// Description: Arithmetic right shift
// =============================================================================

class tc_1_1_8_sra_seq extends uvm_sequence #(rv32i_transaction);
    
    `uvm_object_utils(tc_1_1_8_sra_seq)
    
    function new(string name = "tc_1_1_8_sra_seq");
        super.new(name);
    endfunction
    
    task body();
        rv32i_transaction tr;
        
        `uvm_info(get_type_name(), "Starting SRA sequence", UVM_MEDIUM)
        
        // ======================================================================
        // Test Case: SRA - Arithmetic right shift
        // ======================================================================
        tr = rv32i_transaction::type_id::create("sra_test");
        start_item(tr);
        
        tr.test_name = "SRA Test";
        // TODO: Configure instruction encoding and test values
        // tr.opcode = ...;
        // tr.funct3 = ...;
        // tr.rd = ...;
        // tr.rs1 = ...;
        // tr.rs2 = ...;
        // tr.instruction = {tr.funct7, tr.rs2, tr.rs1, tr.funct3, tr.rd, tr.opcode};
        
        finish_item(tr);
        `uvm_info(get_type_name(), "Sent: SRA test transaction", UVM_HIGH)
        
        `uvm_info(get_type_name(), "SRA sequence completed", UVM_MEDIUM)
        
    endtask

endclass : tc_1_1_8_sra_seq
