// =============================================================================
// Sequence: TC 1.3.1 - LW Instruction
// =============================================================================
// Category: ISA Coverage
// Priority: CRITICAL
// Description: Load word
// =============================================================================

class tc_1_3_1_lw_seq extends uvm_sequence #(rv32i_transaction);
    
    `uvm_object_utils(tc_1_3_1_lw_seq)
    
    function new(string name = "tc_1_3_1_lw_seq");
        super.new(name);
    endfunction
    
    task body();
        rv32i_transaction tr;
        
        `uvm_info(get_type_name(), "Starting LW sequence", UVM_MEDIUM)
        
        // ======================================================================
        // Test Case: LW - Load word
        // ======================================================================
        tr = rv32i_transaction::type_id::create("lw_test");
        start_item(tr);
        
        tr.test_name = "LW Test";
        // TODO: Configure instruction encoding and test values
        // tr.opcode = ...;
        // tr.funct3 = ...;
        // tr.rd = ...;
        // tr.rs1 = ...;
        // tr.rs2 = ...;
        // tr.instruction = {tr.funct7, tr.rs2, tr.rs1, tr.funct3, tr.rd, tr.opcode};
        
        finish_item(tr);
        `uvm_info(get_type_name(), "Sent: LW test transaction", UVM_HIGH)
        
        `uvm_info(get_type_name(), "LW sequence completed", UVM_MEDIUM)
        
    endtask

endclass : tc_1_3_1_lw_seq
