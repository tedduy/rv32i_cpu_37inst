// =============================================================================
// Sequence: TC 4.2.3 - X0_BOTH Instruction
// =============================================================================
// Category: Edge Cases
// Priority: HIGH
// Description: x0 as source and dest
// =============================================================================

class tc_4_2_3_x0_both_seq extends uvm_sequence #(rv32i_transaction);
    
    `uvm_object_utils(tc_4_2_3_x0_both_seq)
    
    function new(string name = "tc_4_2_3_x0_both_seq");
        super.new(name);
    endfunction
    
    task body();
        rv32i_transaction tr;
        
        `uvm_info(get_type_name(), "Starting X0_BOTH sequence", UVM_MEDIUM)
        
        // ======================================================================
        // Test Case: X0_BOTH - x0 as source and dest
        // ======================================================================
        tr = rv32i_transaction::type_id::create("x0_both_test");
        start_item(tr);
        
        tr.test_name = "X0_BOTH Test";
        // TODO: Configure instruction encoding and test values
        // tr.opcode = ...;
        // tr.funct3 = ...;
        // tr.rd = ...;
        // tr.rs1 = ...;
        // tr.rs2 = ...;
        // tr.instruction = {tr.funct7, tr.rs2, tr.rs1, tr.funct3, tr.rd, tr.opcode};
        
        finish_item(tr);
        `uvm_info(get_type_name(), "Sent: X0_BOTH test transaction", UVM_HIGH)
        
        `uvm_info(get_type_name(), "X0_BOTH sequence completed", UVM_MEDIUM)
        
    endtask

endclass : tc_4_2_3_x0_both_seq
